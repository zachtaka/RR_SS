// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: RR_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-08-11 on Sun Jun 17 14:13:58 2018
//=============================================================================
// Description: Package for agent RR
//=============================================================================

package RR_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  `include "RR_trans.sv"
  `include "RR_config.sv"
  `include "RR_driver_wb_fl.sv"
  `include "RR_driver.sv"
  `include "RR_monitor.sv"
  `include "RR_sequencer.sv"
  `include "RR_coverage.sv"
  `include "RR_agent.sv"
  `include "RR_seq_lib.sv"

endpackage : RR_pkg
